//ALU Top Moudle
module alu_top();
endmodule
